// Copyright 2023 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

package riscv_instr_branch;
  localparam logic [31:0] BEQ                = 32'b?????????????????000?????1100011;
  localparam logic [31:0] BNE                = 32'b?????????????????001?????1100011;
  localparam logic [31:0] BLT                = 32'b?????????????????100?????1100011;
  localparam logic [31:0] BGE                = 32'b?????????????????101?????1100011;
  localparam logic [31:0] BLTU               = 32'b?????????????????110?????1100011;
  localparam logic [31:0] BGEU               = 32'b?????????????????111?????1100011;
  localparam logic [31:0] JAL                = 32'b?????????????????????????1101111;
endpackage
